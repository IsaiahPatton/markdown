module markdown

const (
	nl = '\n'
)

pub fn to_plain(input string) string {
	// TODO: markdown to plain text
	mut s := 'todo'
	return s
}
