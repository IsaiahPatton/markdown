module parsers

/**
 * TODO
 */
pub fn parse_referencelink(text string) string {
	mut s := text
	return s
}