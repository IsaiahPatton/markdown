module parsers

/**
 * TODO
 */
pub fn parse_lists(text string) string {
	mut s := text
	return s
}