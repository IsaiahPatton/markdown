module parsers

/**
 * TODO
 */
pub fn parse_italic(text string) string {
	mut s := text
	return s
}