module parsers

/**
 * TODO
 */
pub fn parse_bold(text string) string {
	mut s := text
	return s
}