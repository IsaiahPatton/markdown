module parsers

/**
 * TODO
 */
pub fn parse_blockquote(text string) string {
	mut s := text
	return s
}