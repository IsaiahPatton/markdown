module parsers

/**
 * TODO
 */
pub fn parse_hr(text string) string {
	mut s := text
	return s
}