module parsers

/**
 * TODO
 */
pub fn parse_codeblock(text string) string {
	mut s := text
	return s
}